.title KiCad schematic
.include "C:/AE/MAX16823/_models/C2012C0G1H153J085AA_p.mod"
.include "C:/AE/MAX16823/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/MAX16823/_models/C3216X7R1H105K160AB_p.mod"
.include "C:/AE/MAX16823/_models/MJD31C.spice.txt"
.include "C:/AE/MAX16823/_models/SML-Z14F4T.lib"
.include "C:/AE/MAX16823/_models/SML-Z14U4T.lib"
.include "C:/AE/MAX16823/_models/SML-Z14Y4T.lib"
.include "C:/AE/MAX16823/_models/max16823.lib"
XU8 VCC 0 C3216X7R1H105K160AB_p
V2 /DIMM 0 PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE})
XU1 /REG 0 C2012X7R2A104K125AA_p
XU2 VCC 0 C2012X7R2A104K125AA_p
D9 /Y_3 /SENSE3 SML-Z14Y4T
D8 /Y_2 /Y_3 SML-Z14Y4T
XU7 /Y_1 0 C3216X7R1H105K160AB_p
D5 /Y_1 /Y_2 SML-Z14Y4T
R7 /SENSE3 0 {RSENSE}
R5 /SENSE2 0 {RSENSE}
D6 /R_2 /R_3 SML-Z14U4T
D7 /R_3 /SENSE2 SML-Z14U4T
D3 /R_1 /R_2 SML-Z14U4T
R6 /CHN3 0 {RPD}
Q2 VCC /CHN2 /R_1 MJD31C
Q3 VCC /CHN3 /Y_1 MJD31C
R2 /CHN1 0 {RPD}
R4 /CHN2 0 {RPD}
Q1 VCC /CHN1 /G_1 MJD31C
R3 /SENSE1 0 {RSENSE}
V1 VCC 0 {VSOURCE}
R1 /REG /LEDGOOD {RLG}
XU4 /LGC 0 C2012C0G1H153J085AA_p
XU3 /DIMM /DIMM /DIMM /LEDGOOD VCC /LGC /REG 0 /SENSE3 /SENSE2 /SENSE1 /CHN3 /CHN2 /CHN1 MAX16823
XU6 /R_1 0 C3216X7R1H105K160AB_p
D1 /G_1 /G_2 SML-Z14F4T
D2 /G_2 /G_3 SML-Z14F4T
D4 /G_3 /SENSE1 SML-Z14F4T
XU5 /G_1 0 C3216X7R1H105K160AB_p
.end
